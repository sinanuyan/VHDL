library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity tb_i2c_master is
end tb_i2c_master;

architecture TB of tb_i2c_master is
begin
end TB;