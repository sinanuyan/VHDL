library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity i2c_master is
    port(
        clk: in  std_logic;
        rst_pi : in std_logic
    );
end i2c_master;

architecture rtl of i2c_master is
begin
end rtl;